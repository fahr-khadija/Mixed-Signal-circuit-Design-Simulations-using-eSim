* /home/khadija.fahr/Desktop/mixed_signal/Fahr_clk-RVMyth-Dac/Fahr_clk-RVMyth-Dac.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon 07 Mar 2022 05:03:39 PM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  clk Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ adc_bridge_2		
U5  Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ Net-_U5-Pad5_ Net-_U5-Pad6_ Net-_U5-Pad7_ Net-_U5-Pad8_ Net-_U5-Pad9_ Net-_U5-Pad10_ Net-_U5-Pad11_ Net-_U5-Pad12_ Net-_U5-Pad13_ Net-_U5-Pad14_ Net-_U5-Pad15_ Net-_U5-Pad16_ dac_bridge_8		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ dac_bridge_2		
X2  Net-_U4-Pad4_ Net-_U4-Pad3_ Net-_U5-Pad16_ Net-_U5-Pad15_ Net-_U5-Pad14_ Net-_U5-Pad13_ Net-_U5-Pad12_ Net-_U5-Pad11_ Net-_U5-Pad10_ Net-_U5-Pad9_ out 10bitDAC		
X1  Net-_R1-Pad2_ Net-_R1-Pad1_ c_out clk Clock_pulse_generator		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 1k		
R2  c_out Net-_R1-Pad1_ 10k		
C1  c_out GND 0.1u		
v1  Net-_R1-Pad2_ GND DC		
v2  Net-_U3-Pad2_ GND DC		
u1  c_out plot_v1		
U6  out plot_v1		
U2  clk plot_v1		
U7  Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ Net-_U5-Pad5_ Net-_U5-Pad6_ Net-_U5-Pad7_ Net-_U5-Pad8_ Net-_U4-Pad1_ Net-_U4-Pad2_ fahr_rvmyth		

.end
